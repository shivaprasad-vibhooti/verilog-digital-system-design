module add(input [3:0] A, B,
           output [7:0] result);

    assign result = A + B;

endmodule
